// Sequence class

class seq extends uvm_sequence #(seq_item);
    // task
endclass : seq