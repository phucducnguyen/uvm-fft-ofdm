// Sequence_item class

class seq_item extends uvm_sequence_item;
    rand reg[7:0] rand_seq_item;
    // function new(string name = "seq_item");
    //     super.new(name);
    // endfunction
endclass : seq_item