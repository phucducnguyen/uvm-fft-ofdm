// Sequence_item class

class ifft_seq_item extends uvm_sequence_item;
    
    


endclass : ifft_seq_item