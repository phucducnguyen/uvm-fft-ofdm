// Sequence_item class

class seq_item extends uvm_sequence_item;
    rand reg[7:0] rand_seq_item;
endclass : seq_item